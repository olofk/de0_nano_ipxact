//FIXME: Used to deflatten IRQ bus
module mor1kx_irq
  (input  	 irq0,
   input 	 irq1,
   input 	 irq2,
   input 	 irq3,
   input 	 irq4,
   input 	 irq5,
   input 	 irq6,
   input 	 irq7,
   input 	 irq8,
   input 	 irq9,
   input 	 irq10,
   input 	 irq11,
   input 	 irq12,
   input 	 irq13,
   input 	 irq14,
   input 	 irq15,
   input 	 irq16,
   input 	 irq17,
   input 	 irq18,
   input 	 irq19,
   input 	 irq20,
   input 	 irq21,
   input 	 irq22,
   input 	 irq23,
   input 	 irq24,
   input 	 irq25,
   input 	 irq26,
   input 	 irq27,
   input 	 irq28,
   input 	 irq29,
   input 	 irq30,
   input 	 irq31,

   output [31:0] irq_o);
   
   assign irq_o = {irq31,irq30,irq29,irq28,
		   irq27,irq26,irq25,irq24,
		   irq23,irq22,irq21,irq20,
		   irq19,irq18,irq17,irq16,
		   irq15,irq14,irq13,irq12,
		   irq11,irq10,irq9 ,irq8,
		   irq7 ,irq6 ,irq5 ,irq4,
		   irq3 ,irq2 ,irq1 ,irq0};
endmodule
